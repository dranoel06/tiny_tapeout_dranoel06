module tt_um_dranoel06_SAP1 (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

assign uio_out = 8'b0;   
assign uio_oe  = 8'b0;   


wire ena_unused = ena;
wire [2:0] uio_un_unused = uio_in[6:4];


cpu cpu0(
    .clk(clk),
    .reset(~rst_n),
    .programm_input(ui_in),
    .output_register(uo_out),
    .prog(uio_in[7]),
    .addr(uio_in[3:0])
);


endmodule



